`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.02.2024 16:36:04
// Design Name: 
// Module Name: jump_branch_mod
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module jump_branch_mod(
    input [2:0] func3,
    input [20:0] imm,
    input [63:0] data_rs1,
    input [63:0] data_rs2,
    input [6:0] opcode,
    output [5:0] jump
    );
endmodule
